`include "uvm_macros.svh"

import uvm_pkg::*;

`include "test.sv"

module top;
  initial 
    run_test();




endmodule
