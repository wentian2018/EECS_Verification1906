`ifndef ROUTER_IO__SV
`define ROUTER_IO__SV

interface router_io(input bit clk);

   logic  reset_n ;
   logic [15:0] frame_n ;
   logic [15:0] valid_n ;
   logic [15:0] din ;
   logic [15:0] dout ;
   logic [15:0] busy_n ;
   logic [15:0] valido_n ;
   logic [15:0] frameo_n ;
/*
  Declare a clocking block driven by posedge of signal clock     //
  Add all signals required to connected test program to the DUT  //
  All direction must be with respected to test program           //
*/
   clocking drvClk @(posedge clk);
      output  reset_n;
      output  frame_n;
      output  valid_n;
      output  din;
      input   busy_n;
   endclocking: drvClk

   clocking iMonClk @(posedge clk);
/*
   Add input and output skew in clocking block(optional)
*/
      input  frame_n;
      input  valid_n;
      input  din;
      input  busy_n;
   endclocking: iMonClk

   clocking oMonClk @(posedge clk);
      input  dout;
      input  valido_n;
      input  frameo_n;
   endclocking: oMonClk
/*
   Create modport to connect to test program
   Arguments should list clocking block and all other async signals
*/
   modport driver(clocking drvClk, output reset_n);
   modport imon(clocking iMonClk);
   modport omon(clocking oMonClk);
   modport dut(input clk, reset_n, frame_n, valid_n, din, output dout, busy_n, valido_n, frameo_n);

endinterface: router_io

`endif
